module fe_top 
  #(parameter 
  )
  ( input logic clk_i
  ):



endmodule // fe_top