module priority_encoder
  #( els_p    = -1
    ,width_p  = $clog2(els_p)
  )
  (input  logic [els_p-1:0]           i
  ,output logic [$clog2(els_p)-1:0]   addr_o
  ,output logic                       v_o
  );

  always_comb begin
    v_o     = 1'b0;
    addr_o  = '0;

    for(int unsigned j = 0; j < els_p; j++) begin
      if(i[j]) begin 
        v_o     = 1'b1;
        addr_o  = j;
        break;
      end
    end
  end // always_comb

endmodule // priority_encoder_32

// casez(i)
//       32'b00000000000000000000000000000000: v = 1'b0;
//       32'b???????????????????????????????1: o = 5'd0;
//       32'b??????????????????????????????10: o = 5'd1;
//       32'b?????????????????????????????100: o = 5'd2;
//       32'b????????????????????????????1000: o = 5'd3;
//       32'b???????????????????????????10000: o = 5'd4;
//       32'b??????????????????????????100000: o = 5'd5;
//       32'b?????????????????????????1000000: o = 5'd6;
//       32'b????????????????????????10000000: o = 5'd7;
//       32'b???????????????????????100000000: o = 5'd8;
//       32'b??????????????????????1000000000: o = 5'd9;
//       32'b?????????????????????10000000000: o = 5'd10;
//       32'b????????????????????100000000000: o = 5'd11;
//       32'b???????????????????1000000000000: o = 5'd12;
//       32'b??????????????????10000000000000: o = 5'd13;
//       32'b?????????????????100000000000000: o = 5'd14;
//       32'b????????????????1000000000000000: o = 5'd15;
//       32'b???????????????10000000000000000: o = 5'd16;
//       32'b??????????????100000000000000000: o = 5'd17;
//       32'b?????????????1000000000000000000: o = 5'd18;
//       32'b????????????10000000000000000000: o = 5'd19;
//       32'b???????????100000000000000000000: o = 5'd20;
//       32'b??????????1000000000000000000000: o = 5'd21;
//       32'b?????????10000000000000000000000: o = 5'd22;
//       32'b????????100000000000000000000000: o = 5'd23;
//       32'b???????1000000000000000000000000: o = 5'd24;
//       32'b??????10000000000000000000000000: o = 5'd25;
//       32'b?????100000000000000000000000000: o = 5'd26;
//       32'b????1000000000000000000000000000: o = 5'd27;
//       32'b???10000000000000000000000000000: o = 5'd28;
//       32'b??100000000000000000000000000000: o = 5'd29;
//       32'b?1000000000000000000000000000000: o = 5'd30;
//       32'b10000000000000000000000000000000: o = 5'd31;


// casez(i)
//       16'b0000000000000000: v = 1'b0;
//       16'b???????????????1: o = 5'd0;
//       16'b??????????????10: o = 5'd1;
//       16'b?????????????100: o = 5'd2;
//       16'b????????????1000: o = 5'd3;
//       16'b???????????10000: o = 5'd4;
//       16'b??????????100000: o = 5'd5;
//       16'b?????????1000000: o = 5'd6;
//       16'b????????10000000: o = 5'd7;
//       16'b???????100000000: o = 5'd8;
//       16'b??????1000000000: o = 5'd9;
//       16'b?????10000000000: o = 5'd10;
//       16'b????100000000000: o = 5'd11;
//       16'b???1000000000000: o = 5'd12;
//       16'b??10000000000000: o = 5'd13;
//       16'b?100000000000000: o = 5'd14;
//       16'b1000000000000000: o = 5'd15;

