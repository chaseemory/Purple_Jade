`include "Purple_Jade_pkg.svh"
`include ""

module execute_stage
(input                                      clk_i
 , input                                    reset_i
);
endmodule // execute_stage