module fe_top #(
  )
  (
  ):



endmodule // fe_top