module fe_top 
  #(parameter place_holder = -1
  )
  ( input logic clk_i
  , 
  ):



endmodule // fe_top