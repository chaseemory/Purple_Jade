// A ROM for instructions
// Async Reads
`ifdef VERILATOR
`include "Purple_Jade_pkg.svh"
`endif

module i_rom
  #(localparam  ADDR_WIDTH_LP = $clog2(I_ROM_DEPTH_P)
  )
  ( input   logic [ADDR_WIDTH_LP-1:0] r_addr_i
  , output  logic [WORD_SIZE_P-1:0]   data_o
  );

  logic [WORD_SIZE_P-1:0] mem [I_ROM_DEPTH_P-1:0];

  initial begin
    $readmemb(`TEST_BIN, mem);
  end // initial

  assign data_o = mem[r_addr_i];

endmodule // i_rom