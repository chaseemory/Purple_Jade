`ifndef _ROB_DEF_SVH_
`define _ROB_DEF_SVH_

`include "../common/Purple_Jade_pkg.svh";

`endif